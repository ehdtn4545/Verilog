module incoder(
input d_in;
output d_out;
);


endmodule
