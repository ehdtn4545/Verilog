module decoder(
input d_in;
output d_out;
);

endmodule
